class transaction;
  rand bit a;
  rand bit b;
  rand bit c;
      
    bit sum;
    bit carry;
  
